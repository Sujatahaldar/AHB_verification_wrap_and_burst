`include"AHB_intf.sv"
`include"AHB_TX.sv"
`include"AHB_confg.sv"
`include"AHB_gen.sv"
`include"AHB_drv.sv"
`include"AHB_mon.sv"
`include"AHB_scb.sv"
`include"AHB_cov.sv"
`include "AHB_env.sv"
`include"AHB_tb_top.sv"
`include"AHB_tb.sv"